-- AND gate example for parser tests
entity AND_GATE is
  port (
    A : in  std_logic;
    B : in  std_logic;
    Y : out std_logic
  );
end entity AND_GATE;
