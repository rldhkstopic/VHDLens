-- 마이크로 테스트: entity + port 만
entity AND_GATE is
  port (
    A : in  std_logic;
    B : in  std_logic;
    Y : out std_logic
  );
end entity AND_GATE;
